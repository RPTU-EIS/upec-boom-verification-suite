module tag_array_ext( // @[:anonymous source@96.2]
  input  [5:0]  RW0_addr, // @[:anonymous source@97.4]
  input         RW0_clk, // @[:anonymous source@98.4]
  input  [87:0] RW0_wdata, // @[:anonymous source@99.4]
  output [87:0] RW0_rdata, // @[:anonymous source@100.4]
  input         RW0_en, // @[:anonymous source@101.4]
  input         RW0_wmode, // @[:anonymous source@102.4]
  input  [3:0]  RW0_wmask // @[:anonymous source@103.4]
);
  wire [5:0] mem_0_0_RW0_addr; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@105.4]
  wire [21:0] mem_0_0_RW0_wdata; // @[:anonymous source@105.4]
  wire [21:0] mem_0_0_RW0_rdata; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_wmask; // @[:anonymous source@105.4]
  wire [5:0] mem_0_1_RW0_addr; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_clk; // @[:anonymous source@106.4]
  wire [21:0] mem_0_1_RW0_wdata; // @[:anonymous source@106.4]
  wire [21:0] mem_0_1_RW0_rdata; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_en; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_wmode; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_wmask; // @[:anonymous source@106.4]
  wire [5:0] mem_0_2_RW0_addr; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_clk; // @[:anonymous source@107.4]
  wire [21:0] mem_0_2_RW0_wdata; // @[:anonymous source@107.4]
  wire [21:0] mem_0_2_RW0_rdata; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_en; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_wmode; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_wmask; // @[:anonymous source@107.4]
  wire [5:0] mem_0_3_RW0_addr; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_clk; // @[:anonymous source@108.4]
  wire [21:0] mem_0_3_RW0_wdata; // @[:anonymous source@108.4]
  wire [21:0] mem_0_3_RW0_rdata; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_en; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_wmode; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_wmask; // @[:anonymous source@108.4]
  wire [21:0] RW0_rdata_0_0; // @[:anonymous source@111.4]
  wire [21:0] RW0_rdata_0_1; // @[:anonymous source@118.4]
  wire [21:0] RW0_rdata_0_2; // @[:anonymous source@125.4]
  wire [21:0] RW0_rdata_0_3; // @[:anonymous source@132.4]
  wire [43:0] _GEN_0; // @[:anonymous source@137.4]
  wire [65:0] _GEN_1; // @[:anonymous source@137.4]
  wire [87:0] RW0_rdata_0; // @[:anonymous source@137.4]
  wire [43:0] _GEN_2; // @[:anonymous source@138.4]
  wire [65:0] _GEN_3; // @[:anonymous source@138.4]
  split_tag_array_ext mem_0_0 ( // @[:anonymous source@105.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_tag_array_ext mem_0_1 ( // @[:anonymous source@106.4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_tag_array_ext mem_0_2 ( // @[:anonymous source@107.4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_tag_array_ext mem_0_3 ( // @[:anonymous source@108.4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@111.4]
  assign RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[:anonymous source@118.4]
  assign RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[:anonymous source@125.4]
  assign RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[:anonymous source@132.4]
  assign _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@137.4]
  assign _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@137.4]
  assign RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@137.4]
  assign _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@138.4]
  assign _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@138.4]
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1}; // @[:anonymous source@138.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@110.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@109.4]
  assign mem_0_0_RW0_wdata = RW0_wdata[21:0]; // @[:anonymous source@112.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@115.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@114.4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[:anonymous source@113.4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[:anonymous source@117.4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[:anonymous source@116.4]
  assign mem_0_1_RW0_wdata = RW0_wdata[43:22]; // @[:anonymous source@119.4]
  assign mem_0_1_RW0_en = RW0_en; // @[:anonymous source@122.4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[:anonymous source@121.4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[:anonymous source@120.4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[:anonymous source@124.4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[:anonymous source@123.4]
  assign mem_0_2_RW0_wdata = RW0_wdata[65:44]; // @[:anonymous source@126.4]
  assign mem_0_2_RW0_en = RW0_en; // @[:anonymous source@129.4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[:anonymous source@128.4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[:anonymous source@127.4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[:anonymous source@131.4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[:anonymous source@130.4]
  assign mem_0_3_RW0_wdata = RW0_wdata[87:66]; // @[:anonymous source@133.4]
  assign mem_0_3_RW0_en = RW0_en; // @[:anonymous source@136.4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[:anonymous source@135.4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[:anonymous source@134.4]
endmodule
module array_0_0_ext( // @[:anonymous source@140.2]
  input  [8:0]  W0_addr, // @[:anonymous source@141.4]
  input         W0_clk, // @[:anonymous source@142.4]
  input  [63:0] W0_data, // @[:anonymous source@143.4]
  input         W0_en, // @[:anonymous source@144.4]
  input         W0_mask, // @[:anonymous source@145.4]
  input  [8:0]  R0_addr, // @[:anonymous source@146.4]
  input         R0_clk, // @[:anonymous source@147.4]
  output [63:0] R0_data, // @[:anonymous source@148.4]
  input         R0_en // @[:anonymous source@149.4]
);
  wire [8:0] mem_0_0_W0_addr; // @[:anonymous source@151.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@151.4]
  wire [63:0] mem_0_0_W0_data; // @[:anonymous source@151.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@151.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@151.4]
  wire [8:0] mem_0_0_R0_addr; // @[:anonymous source@151.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@151.4]
  wire [63:0] mem_0_0_R0_data; // @[:anonymous source@151.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@151.4]
  wire [63:0] R0_data_0_0; // @[:anonymous source@159.4]
  wire [63:0] R0_data_0; // @[:anonymous source@161.4]
  split_array_0_0_ext mem_0_0 ( // @[:anonymous source@151.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@159.4]
  assign R0_data_0 = R0_data_0_0; // @[:anonymous source@161.4]
  assign R0_data = mem_0_0_R0_data; // @[:anonymous source@162.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@153.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@152.4]
  assign mem_0_0_W0_data = W0_data; // @[:anonymous source@154.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@156.4]
  assign mem_0_0_W0_mask = W0_mask; // @[:anonymous source@155.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@158.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@157.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@160.4]
endmodule
module tag_array_0_ext( // @[:anonymous source@164.2]
  input  [5:0]  RW0_addr, // @[:anonymous source@165.4]
  input         RW0_clk, // @[:anonymous source@166.4]
  input  [79:0] RW0_wdata, // @[:anonymous source@167.4]
  output [79:0] RW0_rdata, // @[:anonymous source@168.4]
  input         RW0_en, // @[:anonymous source@169.4]
  input         RW0_wmode, // @[:anonymous source@170.4]
  input  [3:0]  RW0_wmask // @[:anonymous source@171.4]
);
  wire [5:0] mem_0_0_RW0_addr; // @[:anonymous source@173.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@173.4]
  wire [19:0] mem_0_0_RW0_wdata; // @[:anonymous source@173.4]
  wire [19:0] mem_0_0_RW0_rdata; // @[:anonymous source@173.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@173.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@173.4]
  wire  mem_0_0_RW0_wmask; // @[:anonymous source@173.4]
  wire [5:0] mem_0_1_RW0_addr; // @[:anonymous source@174.4]
  wire  mem_0_1_RW0_clk; // @[:anonymous source@174.4]
  wire [19:0] mem_0_1_RW0_wdata; // @[:anonymous source@174.4]
  wire [19:0] mem_0_1_RW0_rdata; // @[:anonymous source@174.4]
  wire  mem_0_1_RW0_en; // @[:anonymous source@174.4]
  wire  mem_0_1_RW0_wmode; // @[:anonymous source@174.4]
  wire  mem_0_1_RW0_wmask; // @[:anonymous source@174.4]
  wire [5:0] mem_0_2_RW0_addr; // @[:anonymous source@175.4]
  wire  mem_0_2_RW0_clk; // @[:anonymous source@175.4]
  wire [19:0] mem_0_2_RW0_wdata; // @[:anonymous source@175.4]
  wire [19:0] mem_0_2_RW0_rdata; // @[:anonymous source@175.4]
  wire  mem_0_2_RW0_en; // @[:anonymous source@175.4]
  wire  mem_0_2_RW0_wmode; // @[:anonymous source@175.4]
  wire  mem_0_2_RW0_wmask; // @[:anonymous source@175.4]
  wire [5:0] mem_0_3_RW0_addr; // @[:anonymous source@176.4]
  wire  mem_0_3_RW0_clk; // @[:anonymous source@176.4]
  wire [19:0] mem_0_3_RW0_wdata; // @[:anonymous source@176.4]
  wire [19:0] mem_0_3_RW0_rdata; // @[:anonymous source@176.4]
  wire  mem_0_3_RW0_en; // @[:anonymous source@176.4]
  wire  mem_0_3_RW0_wmode; // @[:anonymous source@176.4]
  wire  mem_0_3_RW0_wmask; // @[:anonymous source@176.4]
  wire [19:0] RW0_rdata_0_0; // @[:anonymous source@179.4]
  wire [19:0] RW0_rdata_0_1; // @[:anonymous source@186.4]
  wire [19:0] RW0_rdata_0_2; // @[:anonymous source@193.4]
  wire [19:0] RW0_rdata_0_3; // @[:anonymous source@200.4]
  wire [39:0] _GEN_0; // @[:anonymous source@205.4]
  wire [59:0] _GEN_1; // @[:anonymous source@205.4]
  wire [79:0] RW0_rdata_0; // @[:anonymous source@205.4]
  wire [39:0] _GEN_2; // @[:anonymous source@206.4]
  wire [59:0] _GEN_3; // @[:anonymous source@206.4]
  split_tag_array_0_ext mem_0_0 ( // @[:anonymous source@173.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_1 ( // @[:anonymous source@174.4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_2 ( // @[:anonymous source@175.4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_3 ( // @[:anonymous source@176.4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@179.4]
  assign RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[:anonymous source@186.4]
  assign RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[:anonymous source@193.4]
  assign RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[:anonymous source@200.4]
  assign _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@205.4]
  assign _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@205.4]
  assign RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@205.4]
  assign _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@206.4]
  assign _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@206.4]
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1}; // @[:anonymous source@206.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@178.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@177.4]
  assign mem_0_0_RW0_wdata = RW0_wdata[19:0]; // @[:anonymous source@180.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@183.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@182.4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[:anonymous source@181.4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[:anonymous source@185.4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[:anonymous source@184.4]
  assign mem_0_1_RW0_wdata = RW0_wdata[39:20]; // @[:anonymous source@187.4]
  assign mem_0_1_RW0_en = RW0_en; // @[:anonymous source@190.4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[:anonymous source@189.4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[:anonymous source@188.4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[:anonymous source@192.4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[:anonymous source@191.4]
  assign mem_0_2_RW0_wdata = RW0_wdata[59:40]; // @[:anonymous source@194.4]
  assign mem_0_2_RW0_en = RW0_en; // @[:anonymous source@197.4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[:anonymous source@196.4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[:anonymous source@195.4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[:anonymous source@199.4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[:anonymous source@198.4]
  assign mem_0_3_RW0_wdata = RW0_wdata[79:60]; // @[:anonymous source@201.4]
  assign mem_0_3_RW0_en = RW0_en; // @[:anonymous source@204.4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[:anonymous source@203.4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[:anonymous source@202.4]
endmodule
module dataArrayWay_0_ext( // @[:anonymous source@208.2]
  input  [8:0]  RW0_addr, // @[:anonymous source@209.4]
  input         RW0_clk, // @[:anonymous source@210.4]
  input  [63:0] RW0_wdata, // @[:anonymous source@211.4]
  output [63:0] RW0_rdata, // @[:anonymous source@212.4]
  input         RW0_en, // @[:anonymous source@213.4]
  input         RW0_wmode // @[:anonymous source@214.4]
);
  wire [8:0] mem_0_0_RW0_addr; // @[:anonymous source@216.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@216.4]
  wire [63:0] mem_0_0_RW0_wdata; // @[:anonymous source@216.4]
  wire [63:0] mem_0_0_RW0_rdata; // @[:anonymous source@216.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@216.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@216.4]
  wire [63:0] RW0_rdata_0_0; // @[:anonymous source@219.4]
  wire [63:0] RW0_rdata_0; // @[:anonymous source@223.4]
  split_dataArrayWay_0_ext mem_0_0 ( // @[:anonymous source@216.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@219.4]
  assign RW0_rdata_0 = RW0_rdata_0_0; // @[:anonymous source@223.4]
  assign RW0_rdata = mem_0_0_RW0_rdata; // @[:anonymous source@224.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@218.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@217.4]
  assign mem_0_0_RW0_wdata = RW0_wdata; // @[:anonymous source@220.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@222.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@221.4]
endmodule
module hi_us_ext( // @[:anonymous source@226.2]
  input  [6:0] W0_addr, // @[:anonymous source@227.4]
  input        W0_clk, // @[:anonymous source@228.4]
  input  [3:0] W0_data, // @[:anonymous source@229.4]
  input        W0_en, // @[:anonymous source@230.4]
  input  [3:0] W0_mask, // @[:anonymous source@231.4]
  input  [6:0] R0_addr, // @[:anonymous source@232.4]
  input        R0_clk, // @[:anonymous source@233.4]
  output [3:0] R0_data, // @[:anonymous source@234.4]
  input        R0_en // @[:anonymous source@235.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@237.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@237.4]
  wire  mem_0_0_W0_data; // @[:anonymous source@237.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@237.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@237.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@237.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@237.4]
  wire  mem_0_0_R0_data; // @[:anonymous source@237.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@237.4]
  wire [6:0] mem_0_1_W0_addr; // @[:anonymous source@238.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@238.4]
  wire  mem_0_1_W0_data; // @[:anonymous source@238.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@238.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@238.4]
  wire [6:0] mem_0_1_R0_addr; // @[:anonymous source@238.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@238.4]
  wire  mem_0_1_R0_data; // @[:anonymous source@238.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@238.4]
  wire [6:0] mem_0_2_W0_addr; // @[:anonymous source@239.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@239.4]
  wire  mem_0_2_W0_data; // @[:anonymous source@239.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@239.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@239.4]
  wire [6:0] mem_0_2_R0_addr; // @[:anonymous source@239.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@239.4]
  wire  mem_0_2_R0_data; // @[:anonymous source@239.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@239.4]
  wire [6:0] mem_0_3_W0_addr; // @[:anonymous source@240.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@240.4]
  wire  mem_0_3_W0_data; // @[:anonymous source@240.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@240.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@240.4]
  wire [6:0] mem_0_3_R0_addr; // @[:anonymous source@240.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@240.4]
  wire  mem_0_3_R0_data; // @[:anonymous source@240.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@240.4]
  wire  R0_data_0_0; // @[:anonymous source@263.4]
  wire  R0_data_0_1; // @[:anonymous source@267.4]
  wire  R0_data_0_2; // @[:anonymous source@271.4]
  wire  R0_data_0_3; // @[:anonymous source@275.4]
  wire [1:0] _GEN_0; // @[:anonymous source@277.4]
  wire [2:0] _GEN_1; // @[:anonymous source@277.4]
  wire [3:0] R0_data_0; // @[:anonymous source@277.4]
  wire [1:0] _GEN_2; // @[:anonymous source@278.4]
  wire [2:0] _GEN_3; // @[:anonymous source@278.4]
  split_hi_us_ext mem_0_0 ( // @[:anonymous source@237.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_hi_us_ext mem_0_1 ( // @[:anonymous source@238.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_hi_us_ext mem_0_2 ( // @[:anonymous source@239.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_hi_us_ext mem_0_3 ( // @[:anonymous source@240.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@263.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@267.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@271.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@275.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@277.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@277.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@277.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@278.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@278.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@278.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@242.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@241.4]
  assign mem_0_0_W0_data = W0_data[0]; // @[:anonymous source@243.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@245.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@244.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@262.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@261.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@264.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@247.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@246.4]
  assign mem_0_1_W0_data = W0_data[1]; // @[:anonymous source@248.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@250.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@249.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@266.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@265.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@268.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@252.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@251.4]
  assign mem_0_2_W0_data = W0_data[2]; // @[:anonymous source@253.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@255.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@254.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@270.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@269.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@272.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@257.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@256.4]
  assign mem_0_3_W0_data = W0_data[3]; // @[:anonymous source@258.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@260.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@259.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@274.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@273.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@276.4]
endmodule
module table_ext( // @[:anonymous source@280.2]
  input  [6:0]  W0_addr, // @[:anonymous source@281.4]
  input         W0_clk, // @[:anonymous source@282.4]
  input  [43:0] W0_data, // @[:anonymous source@283.4]
  input         W0_en, // @[:anonymous source@284.4]
  input  [3:0]  W0_mask, // @[:anonymous source@285.4]
  input  [6:0]  R0_addr, // @[:anonymous source@286.4]
  input         R0_clk, // @[:anonymous source@287.4]
  output [43:0] R0_data, // @[:anonymous source@288.4]
  input         R0_en // @[:anonymous source@289.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@291.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@291.4]
  wire [10:0] mem_0_0_W0_data; // @[:anonymous source@291.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@291.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@291.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@291.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@291.4]
  wire [10:0] mem_0_0_R0_data; // @[:anonymous source@291.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@291.4]
  wire [6:0] mem_0_1_W0_addr; // @[:anonymous source@292.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@292.4]
  wire [10:0] mem_0_1_W0_data; // @[:anonymous source@292.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@292.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@292.4]
  wire [6:0] mem_0_1_R0_addr; // @[:anonymous source@292.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@292.4]
  wire [10:0] mem_0_1_R0_data; // @[:anonymous source@292.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@292.4]
  wire [6:0] mem_0_2_W0_addr; // @[:anonymous source@293.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@293.4]
  wire [10:0] mem_0_2_W0_data; // @[:anonymous source@293.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@293.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@293.4]
  wire [6:0] mem_0_2_R0_addr; // @[:anonymous source@293.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@293.4]
  wire [10:0] mem_0_2_R0_data; // @[:anonymous source@293.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@293.4]
  wire [6:0] mem_0_3_W0_addr; // @[:anonymous source@294.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@294.4]
  wire [10:0] mem_0_3_W0_data; // @[:anonymous source@294.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@294.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@294.4]
  wire [6:0] mem_0_3_R0_addr; // @[:anonymous source@294.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@294.4]
  wire [10:0] mem_0_3_R0_data; // @[:anonymous source@294.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@294.4]
  wire [10:0] R0_data_0_0; // @[:anonymous source@317.4]
  wire [10:0] R0_data_0_1; // @[:anonymous source@321.4]
  wire [10:0] R0_data_0_2; // @[:anonymous source@325.4]
  wire [10:0] R0_data_0_3; // @[:anonymous source@329.4]
  wire [21:0] _GEN_0; // @[:anonymous source@331.4]
  wire [32:0] _GEN_1; // @[:anonymous source@331.4]
  wire [43:0] R0_data_0; // @[:anonymous source@331.4]
  wire [21:0] _GEN_2; // @[:anonymous source@332.4]
  wire [32:0] _GEN_3; // @[:anonymous source@332.4]
  split_table_ext mem_0_0 ( // @[:anonymous source@291.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_table_ext mem_0_1 ( // @[:anonymous source@292.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_table_ext mem_0_2 ( // @[:anonymous source@293.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_table_ext mem_0_3 ( // @[:anonymous source@294.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@317.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@321.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@325.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@329.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@331.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@331.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@331.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@332.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@332.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@332.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@296.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@295.4]
  assign mem_0_0_W0_data = W0_data[10:0]; // @[:anonymous source@297.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@299.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@298.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@316.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@315.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@318.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@301.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@300.4]
  assign mem_0_1_W0_data = W0_data[21:11]; // @[:anonymous source@302.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@304.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@303.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@320.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@319.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@322.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@306.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@305.4]
  assign mem_0_2_W0_data = W0_data[32:22]; // @[:anonymous source@307.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@309.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@308.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@324.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@323.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@326.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@311.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@310.4]
  assign mem_0_3_W0_data = W0_data[43:33]; // @[:anonymous source@312.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@314.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@313.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@328.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@327.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@330.4]
endmodule
module hi_us_0_ext( // @[:anonymous source@334.2]
  input  [7:0] W0_addr, // @[:anonymous source@335.4]
  input        W0_clk, // @[:anonymous source@336.4]
  input  [3:0] W0_data, // @[:anonymous source@337.4]
  input        W0_en, // @[:anonymous source@338.4]
  input  [3:0] W0_mask, // @[:anonymous source@339.4]
  input  [7:0] R0_addr, // @[:anonymous source@340.4]
  input        R0_clk, // @[:anonymous source@341.4]
  output [3:0] R0_data, // @[:anonymous source@342.4]
  input        R0_en // @[:anonymous source@343.4]
);
  wire [7:0] mem_0_0_W0_addr; // @[:anonymous source@345.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@345.4]
  wire  mem_0_0_W0_data; // @[:anonymous source@345.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@345.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@345.4]
  wire [7:0] mem_0_0_R0_addr; // @[:anonymous source@345.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@345.4]
  wire  mem_0_0_R0_data; // @[:anonymous source@345.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@345.4]
  wire [7:0] mem_0_1_W0_addr; // @[:anonymous source@346.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@346.4]
  wire  mem_0_1_W0_data; // @[:anonymous source@346.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@346.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@346.4]
  wire [7:0] mem_0_1_R0_addr; // @[:anonymous source@346.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@346.4]
  wire  mem_0_1_R0_data; // @[:anonymous source@346.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@346.4]
  wire [7:0] mem_0_2_W0_addr; // @[:anonymous source@347.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@347.4]
  wire  mem_0_2_W0_data; // @[:anonymous source@347.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@347.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@347.4]
  wire [7:0] mem_0_2_R0_addr; // @[:anonymous source@347.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@347.4]
  wire  mem_0_2_R0_data; // @[:anonymous source@347.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@347.4]
  wire [7:0] mem_0_3_W0_addr; // @[:anonymous source@348.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@348.4]
  wire  mem_0_3_W0_data; // @[:anonymous source@348.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@348.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@348.4]
  wire [7:0] mem_0_3_R0_addr; // @[:anonymous source@348.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@348.4]
  wire  mem_0_3_R0_data; // @[:anonymous source@348.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@348.4]
  wire  R0_data_0_0; // @[:anonymous source@371.4]
  wire  R0_data_0_1; // @[:anonymous source@375.4]
  wire  R0_data_0_2; // @[:anonymous source@379.4]
  wire  R0_data_0_3; // @[:anonymous source@383.4]
  wire [1:0] _GEN_0; // @[:anonymous source@385.4]
  wire [2:0] _GEN_1; // @[:anonymous source@385.4]
  wire [3:0] R0_data_0; // @[:anonymous source@385.4]
  wire [1:0] _GEN_2; // @[:anonymous source@386.4]
  wire [2:0] _GEN_3; // @[:anonymous source@386.4]
  split_hi_us_0_ext mem_0_0 ( // @[:anonymous source@345.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_hi_us_0_ext mem_0_1 ( // @[:anonymous source@346.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_hi_us_0_ext mem_0_2 ( // @[:anonymous source@347.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_hi_us_0_ext mem_0_3 ( // @[:anonymous source@348.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@371.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@375.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@379.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@383.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@385.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@385.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@385.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@386.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@386.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@386.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@350.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@349.4]
  assign mem_0_0_W0_data = W0_data[0]; // @[:anonymous source@351.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@353.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@352.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@370.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@369.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@372.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@355.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@354.4]
  assign mem_0_1_W0_data = W0_data[1]; // @[:anonymous source@356.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@358.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@357.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@374.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@373.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@376.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@360.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@359.4]
  assign mem_0_2_W0_data = W0_data[2]; // @[:anonymous source@361.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@363.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@362.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@378.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@377.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@380.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@365.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@364.4]
  assign mem_0_3_W0_data = W0_data[3]; // @[:anonymous source@366.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@368.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@367.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@382.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@381.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@384.4]
endmodule
module table_0_ext( // @[:anonymous source@388.2]
  input  [7:0]  W0_addr, // @[:anonymous source@389.4]
  input         W0_clk, // @[:anonymous source@390.4]
  input  [47:0] W0_data, // @[:anonymous source@391.4]
  input         W0_en, // @[:anonymous source@392.4]
  input  [3:0]  W0_mask, // @[:anonymous source@393.4]
  input  [7:0]  R0_addr, // @[:anonymous source@394.4]
  input         R0_clk, // @[:anonymous source@395.4]
  output [47:0] R0_data, // @[:anonymous source@396.4]
  input         R0_en // @[:anonymous source@397.4]
);
  wire [7:0] mem_0_0_W0_addr; // @[:anonymous source@399.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@399.4]
  wire [11:0] mem_0_0_W0_data; // @[:anonymous source@399.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@399.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@399.4]
  wire [7:0] mem_0_0_R0_addr; // @[:anonymous source@399.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@399.4]
  wire [11:0] mem_0_0_R0_data; // @[:anonymous source@399.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@399.4]
  wire [7:0] mem_0_1_W0_addr; // @[:anonymous source@400.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@400.4]
  wire [11:0] mem_0_1_W0_data; // @[:anonymous source@400.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@400.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@400.4]
  wire [7:0] mem_0_1_R0_addr; // @[:anonymous source@400.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@400.4]
  wire [11:0] mem_0_1_R0_data; // @[:anonymous source@400.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@400.4]
  wire [7:0] mem_0_2_W0_addr; // @[:anonymous source@401.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@401.4]
  wire [11:0] mem_0_2_W0_data; // @[:anonymous source@401.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@401.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@401.4]
  wire [7:0] mem_0_2_R0_addr; // @[:anonymous source@401.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@401.4]
  wire [11:0] mem_0_2_R0_data; // @[:anonymous source@401.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@401.4]
  wire [7:0] mem_0_3_W0_addr; // @[:anonymous source@402.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@402.4]
  wire [11:0] mem_0_3_W0_data; // @[:anonymous source@402.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@402.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@402.4]
  wire [7:0] mem_0_3_R0_addr; // @[:anonymous source@402.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@402.4]
  wire [11:0] mem_0_3_R0_data; // @[:anonymous source@402.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@402.4]
  wire [11:0] R0_data_0_0; // @[:anonymous source@425.4]
  wire [11:0] R0_data_0_1; // @[:anonymous source@429.4]
  wire [11:0] R0_data_0_2; // @[:anonymous source@433.4]
  wire [11:0] R0_data_0_3; // @[:anonymous source@437.4]
  wire [23:0] _GEN_0; // @[:anonymous source@439.4]
  wire [35:0] _GEN_1; // @[:anonymous source@439.4]
  wire [47:0] R0_data_0; // @[:anonymous source@439.4]
  wire [23:0] _GEN_2; // @[:anonymous source@440.4]
  wire [35:0] _GEN_3; // @[:anonymous source@440.4]
  split_table_0_ext mem_0_0 ( // @[:anonymous source@399.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_table_0_ext mem_0_1 ( // @[:anonymous source@400.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_table_0_ext mem_0_2 ( // @[:anonymous source@401.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_table_0_ext mem_0_3 ( // @[:anonymous source@402.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@425.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@429.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@433.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@437.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@439.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@439.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@439.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@440.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@440.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@440.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@404.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@403.4]
  assign mem_0_0_W0_data = W0_data[11:0]; // @[:anonymous source@405.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@407.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@406.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@424.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@423.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@426.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@409.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@408.4]
  assign mem_0_1_W0_data = W0_data[23:12]; // @[:anonymous source@410.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@412.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@411.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@428.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@427.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@430.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@414.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@413.4]
  assign mem_0_2_W0_data = W0_data[35:24]; // @[:anonymous source@415.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@417.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@416.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@432.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@431.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@434.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@419.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@418.4]
  assign mem_0_3_W0_data = W0_data[47:36]; // @[:anonymous source@420.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@422.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@421.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@436.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@435.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@438.4]
endmodule
module table_1_ext( // @[:anonymous source@442.2]
  input  [6:0]  W0_addr, // @[:anonymous source@443.4]
  input         W0_clk, // @[:anonymous source@444.4]
  input  [51:0] W0_data, // @[:anonymous source@445.4]
  input         W0_en, // @[:anonymous source@446.4]
  input  [3:0]  W0_mask, // @[:anonymous source@447.4]
  input  [6:0]  R0_addr, // @[:anonymous source@448.4]
  input         R0_clk, // @[:anonymous source@449.4]
  output [51:0] R0_data, // @[:anonymous source@450.4]
  input         R0_en // @[:anonymous source@451.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@453.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@453.4]
  wire [12:0] mem_0_0_W0_data; // @[:anonymous source@453.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@453.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@453.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@453.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@453.4]
  wire [12:0] mem_0_0_R0_data; // @[:anonymous source@453.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@453.4]
  wire [6:0] mem_0_1_W0_addr; // @[:anonymous source@454.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@454.4]
  wire [12:0] mem_0_1_W0_data; // @[:anonymous source@454.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@454.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@454.4]
  wire [6:0] mem_0_1_R0_addr; // @[:anonymous source@454.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@454.4]
  wire [12:0] mem_0_1_R0_data; // @[:anonymous source@454.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@454.4]
  wire [6:0] mem_0_2_W0_addr; // @[:anonymous source@455.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@455.4]
  wire [12:0] mem_0_2_W0_data; // @[:anonymous source@455.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@455.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@455.4]
  wire [6:0] mem_0_2_R0_addr; // @[:anonymous source@455.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@455.4]
  wire [12:0] mem_0_2_R0_data; // @[:anonymous source@455.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@455.4]
  wire [6:0] mem_0_3_W0_addr; // @[:anonymous source@456.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@456.4]
  wire [12:0] mem_0_3_W0_data; // @[:anonymous source@456.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@456.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@456.4]
  wire [6:0] mem_0_3_R0_addr; // @[:anonymous source@456.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@456.4]
  wire [12:0] mem_0_3_R0_data; // @[:anonymous source@456.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@456.4]
  wire [12:0] R0_data_0_0; // @[:anonymous source@479.4]
  wire [12:0] R0_data_0_1; // @[:anonymous source@483.4]
  wire [12:0] R0_data_0_2; // @[:anonymous source@487.4]
  wire [12:0] R0_data_0_3; // @[:anonymous source@491.4]
  wire [25:0] _GEN_0; // @[:anonymous source@493.4]
  wire [38:0] _GEN_1; // @[:anonymous source@493.4]
  wire [51:0] R0_data_0; // @[:anonymous source@493.4]
  wire [25:0] _GEN_2; // @[:anonymous source@494.4]
  wire [38:0] _GEN_3; // @[:anonymous source@494.4]
  split_table_1_ext mem_0_0 ( // @[:anonymous source@453.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_table_1_ext mem_0_1 ( // @[:anonymous source@454.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_table_1_ext mem_0_2 ( // @[:anonymous source@455.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_table_1_ext mem_0_3 ( // @[:anonymous source@456.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@479.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@483.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@487.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@491.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@493.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@493.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@493.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@494.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@494.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@494.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@458.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@457.4]
  assign mem_0_0_W0_data = W0_data[12:0]; // @[:anonymous source@459.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@461.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@460.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@478.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@477.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@480.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@463.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@462.4]
  assign mem_0_1_W0_data = W0_data[25:13]; // @[:anonymous source@464.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@466.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@465.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@482.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@481.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@484.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@468.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@467.4]
  assign mem_0_2_W0_data = W0_data[38:26]; // @[:anonymous source@469.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@471.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@470.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@486.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@485.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@488.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@473.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@472.4]
  assign mem_0_3_W0_data = W0_data[51:39]; // @[:anonymous source@474.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@476.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@475.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@490.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@489.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@492.4]
endmodule
module meta_0_ext( // @[:anonymous source@496.2]
  input  [6:0]   W0_addr, // @[:anonymous source@497.4]
  input          W0_clk, // @[:anonymous source@498.4]
  input  [123:0] W0_data, // @[:anonymous source@499.4]
  input          W0_en, // @[:anonymous source@500.4]
  input  [3:0]   W0_mask, // @[:anonymous source@501.4]
  input  [6:0]   R0_addr, // @[:anonymous source@502.4]
  input          R0_clk, // @[:anonymous source@503.4]
  output [123:0] R0_data, // @[:anonymous source@504.4]
  input          R0_en // @[:anonymous source@505.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@507.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@507.4]
  wire [30:0] mem_0_0_W0_data; // @[:anonymous source@507.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@507.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@507.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@507.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@507.4]
  wire [30:0] mem_0_0_R0_data; // @[:anonymous source@507.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@507.4]
  wire [6:0] mem_0_1_W0_addr; // @[:anonymous source@508.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@508.4]
  wire [30:0] mem_0_1_W0_data; // @[:anonymous source@508.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@508.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@508.4]
  wire [6:0] mem_0_1_R0_addr; // @[:anonymous source@508.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@508.4]
  wire [30:0] mem_0_1_R0_data; // @[:anonymous source@508.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@508.4]
  wire [6:0] mem_0_2_W0_addr; // @[:anonymous source@509.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@509.4]
  wire [30:0] mem_0_2_W0_data; // @[:anonymous source@509.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@509.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@509.4]
  wire [6:0] mem_0_2_R0_addr; // @[:anonymous source@509.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@509.4]
  wire [30:0] mem_0_2_R0_data; // @[:anonymous source@509.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@509.4]
  wire [6:0] mem_0_3_W0_addr; // @[:anonymous source@510.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@510.4]
  wire [30:0] mem_0_3_W0_data; // @[:anonymous source@510.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@510.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@510.4]
  wire [6:0] mem_0_3_R0_addr; // @[:anonymous source@510.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@510.4]
  wire [30:0] mem_0_3_R0_data; // @[:anonymous source@510.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@510.4]
  wire [30:0] R0_data_0_0; // @[:anonymous source@533.4]
  wire [30:0] R0_data_0_1; // @[:anonymous source@537.4]
  wire [30:0] R0_data_0_2; // @[:anonymous source@541.4]
  wire [30:0] R0_data_0_3; // @[:anonymous source@545.4]
  wire [61:0] _GEN_0; // @[:anonymous source@547.4]
  wire [92:0] _GEN_1; // @[:anonymous source@547.4]
  wire [123:0] R0_data_0; // @[:anonymous source@547.4]
  wire [61:0] _GEN_2; // @[:anonymous source@548.4]
  wire [92:0] _GEN_3; // @[:anonymous source@548.4]
  split_meta_0_ext mem_0_0 ( // @[:anonymous source@507.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_meta_0_ext mem_0_1 ( // @[:anonymous source@508.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_meta_0_ext mem_0_2 ( // @[:anonymous source@509.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_meta_0_ext mem_0_3 ( // @[:anonymous source@510.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@533.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@537.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@541.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@545.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@547.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@547.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@547.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@548.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@548.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@548.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@512.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@511.4]
  assign mem_0_0_W0_data = W0_data[30:0]; // @[:anonymous source@513.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@515.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@514.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@532.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@531.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@534.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@517.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@516.4]
  assign mem_0_1_W0_data = W0_data[61:31]; // @[:anonymous source@518.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@520.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@519.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@536.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@535.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@538.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@522.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@521.4]
  assign mem_0_2_W0_data = W0_data[92:62]; // @[:anonymous source@523.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@525.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@524.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@540.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@539.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@542.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@527.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@526.4]
  assign mem_0_3_W0_data = W0_data[123:93]; // @[:anonymous source@528.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@530.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@529.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@544.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@543.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@546.4]
endmodule
module btb_0_ext( // @[:anonymous source@550.2]
  input  [6:0]  W0_addr, // @[:anonymous source@551.4]
  input         W0_clk, // @[:anonymous source@552.4]
  input  [55:0] W0_data, // @[:anonymous source@553.4]
  input         W0_en, // @[:anonymous source@554.4]
  input  [3:0]  W0_mask, // @[:anonymous source@555.4]
  input  [6:0]  R0_addr, // @[:anonymous source@556.4]
  input         R0_clk, // @[:anonymous source@557.4]
  output [55:0] R0_data, // @[:anonymous source@558.4]
  input         R0_en // @[:anonymous source@559.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@561.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@561.4]
  wire [13:0] mem_0_0_W0_data; // @[:anonymous source@561.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@561.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@561.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@561.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@561.4]
  wire [13:0] mem_0_0_R0_data; // @[:anonymous source@561.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@561.4]
  wire [6:0] mem_0_1_W0_addr; // @[:anonymous source@562.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@562.4]
  wire [13:0] mem_0_1_W0_data; // @[:anonymous source@562.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@562.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@562.4]
  wire [6:0] mem_0_1_R0_addr; // @[:anonymous source@562.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@562.4]
  wire [13:0] mem_0_1_R0_data; // @[:anonymous source@562.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@562.4]
  wire [6:0] mem_0_2_W0_addr; // @[:anonymous source@563.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@563.4]
  wire [13:0] mem_0_2_W0_data; // @[:anonymous source@563.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@563.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@563.4]
  wire [6:0] mem_0_2_R0_addr; // @[:anonymous source@563.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@563.4]
  wire [13:0] mem_0_2_R0_data; // @[:anonymous source@563.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@563.4]
  wire [6:0] mem_0_3_W0_addr; // @[:anonymous source@564.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@564.4]
  wire [13:0] mem_0_3_W0_data; // @[:anonymous source@564.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@564.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@564.4]
  wire [6:0] mem_0_3_R0_addr; // @[:anonymous source@564.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@564.4]
  wire [13:0] mem_0_3_R0_data; // @[:anonymous source@564.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@564.4]
  wire [13:0] R0_data_0_0; // @[:anonymous source@587.4]
  wire [13:0] R0_data_0_1; // @[:anonymous source@591.4]
  wire [13:0] R0_data_0_2; // @[:anonymous source@595.4]
  wire [13:0] R0_data_0_3; // @[:anonymous source@599.4]
  wire [27:0] _GEN_0; // @[:anonymous source@601.4]
  wire [41:0] _GEN_1; // @[:anonymous source@601.4]
  wire [55:0] R0_data_0; // @[:anonymous source@601.4]
  wire [27:0] _GEN_2; // @[:anonymous source@602.4]
  wire [41:0] _GEN_3; // @[:anonymous source@602.4]
  split_btb_0_ext mem_0_0 ( // @[:anonymous source@561.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_btb_0_ext mem_0_1 ( // @[:anonymous source@562.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_btb_0_ext mem_0_2 ( // @[:anonymous source@563.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_btb_0_ext mem_0_3 ( // @[:anonymous source@564.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@587.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@591.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@595.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@599.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@601.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@601.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@601.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@602.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@602.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@602.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@566.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@565.4]
  assign mem_0_0_W0_data = W0_data[13:0]; // @[:anonymous source@567.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@569.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@568.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@586.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@585.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@588.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@571.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@570.4]
  assign mem_0_1_W0_data = W0_data[27:14]; // @[:anonymous source@572.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@574.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@573.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@590.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@589.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@592.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@576.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@575.4]
  assign mem_0_2_W0_data = W0_data[41:28]; // @[:anonymous source@577.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@579.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@578.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@594.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@593.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@596.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@581.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@580.4]
  assign mem_0_3_W0_data = W0_data[55:42]; // @[:anonymous source@582.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@584.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@583.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@598.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@597.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@600.4]
endmodule
module ebtb_ext( // @[:anonymous source@604.2]
  input  [6:0]  W0_addr, // @[:anonymous source@605.4]
  input         W0_clk, // @[:anonymous source@606.4]
  input  [39:0] W0_data, // @[:anonymous source@607.4]
  input         W0_en, // @[:anonymous source@608.4]
  input  [6:0]  R0_addr, // @[:anonymous source@609.4]
  input         R0_clk, // @[:anonymous source@610.4]
  output [39:0] R0_data, // @[:anonymous source@611.4]
  input         R0_en // @[:anonymous source@612.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@614.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@614.4]
  wire [39:0] mem_0_0_W0_data; // @[:anonymous source@614.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@614.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@614.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@614.4]
  wire [39:0] mem_0_0_R0_data; // @[:anonymous source@614.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@614.4]
  wire [39:0] R0_data_0_0; // @[:anonymous source@621.4]
  wire [39:0] R0_data_0; // @[:anonymous source@623.4]
  split_ebtb_ext mem_0_0 ( // @[:anonymous source@614.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@621.4]
  assign R0_data_0 = R0_data_0_0; // @[:anonymous source@623.4]
  assign R0_data = mem_0_0_R0_data; // @[:anonymous source@624.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@616.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@615.4]
  assign mem_0_0_W0_data = W0_data; // @[:anonymous source@617.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@618.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@620.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@619.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@622.4]
endmodule
module data_ext( // @[:anonymous source@626.2]
  input  [10:0] W0_addr, // @[:anonymous source@627.4]
  input         W0_clk, // @[:anonymous source@628.4]
  input  [7:0]  W0_data, // @[:anonymous source@629.4]
  input         W0_en, // @[:anonymous source@630.4]
  input  [3:0]  W0_mask, // @[:anonymous source@631.4]
  input  [10:0] R0_addr, // @[:anonymous source@632.4]
  input         R0_clk, // @[:anonymous source@633.4]
  output [7:0]  R0_data, // @[:anonymous source@634.4]
  input         R0_en // @[:anonymous source@635.4]
);
  wire [10:0] mem_0_0_W0_addr; // @[:anonymous source@637.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@637.4]
  wire [1:0] mem_0_0_W0_data; // @[:anonymous source@637.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@637.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@637.4]
  wire [10:0] mem_0_0_R0_addr; // @[:anonymous source@637.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@637.4]
  wire [1:0] mem_0_0_R0_data; // @[:anonymous source@637.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@637.4]
  wire [10:0] mem_0_1_W0_addr; // @[:anonymous source@638.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@638.4]
  wire [1:0] mem_0_1_W0_data; // @[:anonymous source@638.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@638.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@638.4]
  wire [10:0] mem_0_1_R0_addr; // @[:anonymous source@638.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@638.4]
  wire [1:0] mem_0_1_R0_data; // @[:anonymous source@638.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@638.4]
  wire [10:0] mem_0_2_W0_addr; // @[:anonymous source@639.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@639.4]
  wire [1:0] mem_0_2_W0_data; // @[:anonymous source@639.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@639.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@639.4]
  wire [10:0] mem_0_2_R0_addr; // @[:anonymous source@639.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@639.4]
  wire [1:0] mem_0_2_R0_data; // @[:anonymous source@639.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@639.4]
  wire [10:0] mem_0_3_W0_addr; // @[:anonymous source@640.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@640.4]
  wire [1:0] mem_0_3_W0_data; // @[:anonymous source@640.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@640.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@640.4]
  wire [10:0] mem_0_3_R0_addr; // @[:anonymous source@640.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@640.4]
  wire [1:0] mem_0_3_R0_data; // @[:anonymous source@640.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@640.4]
  wire [1:0] R0_data_0_0; // @[:anonymous source@663.4]
  wire [1:0] R0_data_0_1; // @[:anonymous source@667.4]
  wire [1:0] R0_data_0_2; // @[:anonymous source@671.4]
  wire [1:0] R0_data_0_3; // @[:anonymous source@675.4]
  wire [3:0] _GEN_0; // @[:anonymous source@677.4]
  wire [5:0] _GEN_1; // @[:anonymous source@677.4]
  wire [7:0] R0_data_0; // @[:anonymous source@677.4]
  wire [3:0] _GEN_2; // @[:anonymous source@678.4]
  wire [5:0] _GEN_3; // @[:anonymous source@678.4]
  split_data_ext mem_0_0 ( // @[:anonymous source@637.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_data_ext mem_0_1 ( // @[:anonymous source@638.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_data_ext mem_0_2 ( // @[:anonymous source@639.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_data_ext mem_0_3 ( // @[:anonymous source@640.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@663.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@667.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@671.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@675.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@677.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@677.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@677.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@678.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@678.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@678.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@642.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@641.4]
  assign mem_0_0_W0_data = W0_data[1:0]; // @[:anonymous source@643.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@645.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@644.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@662.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@661.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@664.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@647.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@646.4]
  assign mem_0_1_W0_data = W0_data[3:2]; // @[:anonymous source@648.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@650.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@649.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@666.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@665.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@668.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@652.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@651.4]
  assign mem_0_2_W0_data = W0_data[5:4]; // @[:anonymous source@653.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@655.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@654.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@670.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@669.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@672.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@657.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@656.4]
  assign mem_0_3_W0_data = W0_data[7:6]; // @[:anonymous source@658.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@660.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@659.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@674.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@673.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@676.4]
endmodule
module meta_ext( // @[:anonymous source@680.2]
  input  [4:0]   W0_addr, // @[:anonymous source@681.4]
  input          W0_clk, // @[:anonymous source@682.4]
  input  [119:0] W0_data, // @[:anonymous source@683.4]
  input          W0_en, // @[:anonymous source@684.4]
  input  [4:0]   R0_addr, // @[:anonymous source@685.4]
  input          R0_clk, // @[:anonymous source@686.4]
  output [119:0] R0_data, // @[:anonymous source@687.4]
  input          R0_en // @[:anonymous source@688.4]
);
  wire [4:0] mem_0_0_W0_addr; // @[:anonymous source@690.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@690.4]
  wire [119:0] mem_0_0_W0_data; // @[:anonymous source@690.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@690.4]
  wire [4:0] mem_0_0_R0_addr; // @[:anonymous source@690.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@690.4]
  wire [119:0] mem_0_0_R0_data; // @[:anonymous source@690.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@690.4]
  wire [119:0] R0_data_0_0; // @[:anonymous source@697.4]
  wire [119:0] R0_data_0; // @[:anonymous source@699.4]
  split_meta_ext mem_0_0 ( // @[:anonymous source@690.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@697.4]
  assign R0_data_0 = R0_data_0_0; // @[:anonymous source@699.4]
  assign R0_data = mem_0_0_R0_data; // @[:anonymous source@700.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@692.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@691.4]
  assign mem_0_0_W0_data = W0_data; // @[:anonymous source@693.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@694.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@696.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@695.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@698.4]
endmodule
module ghist_0_ext( // @[:anonymous source@702.2]
  input  [4:0]  W0_addr, // @[:anonymous source@703.4]
  input         W0_clk, // @[:anonymous source@704.4]
  input  [71:0] W0_data, // @[:anonymous source@705.4]
  input         W0_en, // @[:anonymous source@706.4]
  input  [4:0]  R0_addr, // @[:anonymous source@707.4]
  input         R0_clk, // @[:anonymous source@708.4]
  output [71:0] R0_data, // @[:anonymous source@709.4]
  input         R0_en // @[:anonymous source@710.4]
);
  wire [4:0] mem_0_0_W0_addr; // @[:anonymous source@712.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@712.4]
  wire [71:0] mem_0_0_W0_data; // @[:anonymous source@712.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@712.4]
  wire [4:0] mem_0_0_R0_addr; // @[:anonymous source@712.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@712.4]
  wire [71:0] mem_0_0_R0_data; // @[:anonymous source@712.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@712.4]
  wire [71:0] R0_data_0_0; // @[:anonymous source@719.4]
  wire [71:0] R0_data_0; // @[:anonymous source@721.4]
  split_ghist_0_ext mem_0_0 ( // @[:anonymous source@712.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@719.4]
  assign R0_data_0 = R0_data_0_0; // @[:anonymous source@721.4]
  assign R0_data = mem_0_0_R0_data; // @[:anonymous source@722.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@714.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@713.4]
  assign mem_0_0_W0_data = W0_data; // @[:anonymous source@715.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@716.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@718.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@717.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@720.4]
endmodule
module rob_debug_inst_mem_ext( // @[:anonymous source@724.2]
  input  [4:0]  W0_addr, // @[:anonymous source@725.4]
  input         W0_clk, // @[:anonymous source@726.4]
  input  [63:0] W0_data, // @[:anonymous source@727.4]
  input         W0_en, // @[:anonymous source@728.4]
  input  [1:0]  W0_mask, // @[:anonymous source@729.4]
  input  [4:0]  R0_addr, // @[:anonymous source@730.4]
  input         R0_clk, // @[:anonymous source@731.4]
  output [63:0] R0_data, // @[:anonymous source@732.4]
  input         R0_en // @[:anonymous source@733.4]
);
  wire [4:0] mem_0_0_W0_addr; // @[:anonymous source@735.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@735.4]
  wire [31:0] mem_0_0_W0_data; // @[:anonymous source@735.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@735.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@735.4]
  wire [4:0] mem_0_0_R0_addr; // @[:anonymous source@735.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@735.4]
  wire [31:0] mem_0_0_R0_data; // @[:anonymous source@735.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@735.4]
  wire [4:0] mem_0_1_W0_addr; // @[:anonymous source@736.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@736.4]
  wire [31:0] mem_0_1_W0_data; // @[:anonymous source@736.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@736.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@736.4]
  wire [4:0] mem_0_1_R0_addr; // @[:anonymous source@736.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@736.4]
  wire [31:0] mem_0_1_R0_data; // @[:anonymous source@736.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@736.4]
  wire [31:0] R0_data_0_0; // @[:anonymous source@749.4]
  wire [31:0] R0_data_0_1; // @[:anonymous source@753.4]
  wire [63:0] R0_data_0; // @[:anonymous source@755.4]
  split_rob_debug_inst_mem_ext mem_0_0 ( // @[:anonymous source@735.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_rob_debug_inst_mem_ext mem_0_1 ( // @[:anonymous source@736.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@749.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@753.4]
  assign R0_data_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@755.4]
  assign R0_data = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@756.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@738.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@737.4]
  assign mem_0_0_W0_data = W0_data[31:0]; // @[:anonymous source@739.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@741.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@740.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@748.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@747.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@750.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@743.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@742.4]
  assign mem_0_1_W0_data = W0_data[63:32]; // @[:anonymous source@744.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@746.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@745.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@752.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@751.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@754.4]
endmodule
module l2_tlb_ram_ext( // @[:anonymous source@758.2]
  input  [9:0]  RW0_addr, // @[:anonymous source@759.4]
  input         RW0_clk, // @[:anonymous source@760.4]
  input  [43:0] RW0_wdata, // @[:anonymous source@761.4]
  output [43:0] RW0_rdata, // @[:anonymous source@762.4]
  input         RW0_en, // @[:anonymous source@763.4]
  input         RW0_wmode // @[:anonymous source@764.4]
);
  wire [9:0] mem_0_0_RW0_addr; // @[:anonymous source@766.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@766.4]
  wire [43:0] mem_0_0_RW0_wdata; // @[:anonymous source@766.4]
  wire [43:0] mem_0_0_RW0_rdata; // @[:anonymous source@766.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@766.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@766.4]
  wire [43:0] RW0_rdata_0_0; // @[:anonymous source@769.4]
  wire [43:0] RW0_rdata_0; // @[:anonymous source@773.4]
  split_l2_tlb_ram_ext mem_0_0 ( // @[:anonymous source@766.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@769.4]
  assign RW0_rdata_0 = RW0_rdata_0_0; // @[:anonymous source@773.4]
  assign RW0_rdata = mem_0_0_RW0_rdata; // @[:anonymous source@774.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@768.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@767.4]
  assign mem_0_0_RW0_wdata = RW0_wdata; // @[:anonymous source@770.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@772.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@771.4]
endmodule
module split_tag_array_ext( // @[:anonymous source@823.2]
  input  [5:0]  RW0_addr, // @[:anonymous source@824.4]
  input         RW0_clk, // @[:anonymous source@825.4]
  input  [21:0] RW0_wdata, // @[:anonymous source@826.4]
  output [21:0] RW0_rdata, // @[:anonymous source@827.4]
  input         RW0_en, // @[:anonymous source@828.4]
  input         RW0_wmode, // @[:anonymous source@829.4]
  input         RW0_wmask // @[:anonymous source@830.4]
);
  reg [21:0] ram [0:63]; // @[:anonymous source@832.4]
  reg [31:0] _RAND_0;
  wire [21:0] ram_RW_0_r_data; // @[:anonymous source@832.4]
  wire [5:0] ram_RW_0_r_addr; // @[:anonymous source@832.4]
  wire [21:0] ram_RW_0_w_data; // @[:anonymous source@832.4]
  wire [5:0] ram_RW_0_w_addr; // @[:anonymous source@832.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@832.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@832.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [5:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@832.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@844.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@832.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_array_0_0_ext( // @[:anonymous source@847.2]
  input  [8:0]  W0_addr, // @[:anonymous source@848.4]
  input         W0_clk, // @[:anonymous source@849.4]
  input  [63:0] W0_data, // @[:anonymous source@850.4]
  input         W0_en, // @[:anonymous source@851.4]
  input         W0_mask, // @[:anonymous source@852.4]
  input  [8:0]  R0_addr, // @[:anonymous source@853.4]
  input         R0_clk, // @[:anonymous source@854.4]
  output [63:0] R0_data, // @[:anonymous source@855.4]
  input         R0_en // @[:anonymous source@856.4]
);
  reg [63:0] ram [0:63]; // @[:anonymous source@858.4]
  reg [63:0] _RAND_0;
  wire [63:0] ram_R_0_data; // @[:anonymous source@858.4]
  wire [8:0] ram_R_0_addr; // @[:anonymous source@858.4]
  wire [63:0] ram_W_0_data; // @[:anonymous source@858.4]
  wire [8:0] ram_W_0_addr; // @[:anonymous source@858.4]
  wire  ram_W_0_mask; // @[:anonymous source@858.4]
  wire  ram_W_0_en; // @[:anonymous source@858.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [8:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@858.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@869.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@858.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_tag_array_0_ext( // @[:anonymous source@876.2]
  input  [5:0]  RW0_addr, // @[:anonymous source@877.4]
  input         RW0_clk, // @[:anonymous source@878.4]
  input  [19:0] RW0_wdata, // @[:anonymous source@879.4]
  output [19:0] RW0_rdata, // @[:anonymous source@880.4]
  input         RW0_en, // @[:anonymous source@881.4]
  input         RW0_wmode, // @[:anonymous source@882.4]
  input         RW0_wmask // @[:anonymous source@883.4]
);
  reg [19:0] ram [0:63]; // @[:anonymous source@885.4]
  reg [31:0] _RAND_0;
  wire [19:0] ram_RW_0_r_data; // @[:anonymous source@885.4]
  wire [5:0] ram_RW_0_r_addr; // @[:anonymous source@885.4]
  wire [19:0] ram_RW_0_w_data; // @[:anonymous source@885.4]
  wire [5:0] ram_RW_0_w_addr; // @[:anonymous source@885.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@885.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@885.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [5:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@885.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@897.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[19:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@885.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_dataArrayWay_0_ext( // @[:anonymous source@900.2]
  input  [8:0]  RW0_addr, // @[:anonymous source@901.4]
  input         RW0_clk, // @[:anonymous source@902.4]
  input  [63:0] RW0_wdata, // @[:anonymous source@903.4]
  output [63:0] RW0_rdata, // @[:anonymous source@904.4]
  input         RW0_en, // @[:anonymous source@905.4]
  input         RW0_wmode // @[:anonymous source@906.4]
);
  reg [63:0] ram [0:63]; // @[:anonymous source@908.4]
  reg [63:0] _RAND_0;
  wire [63:0] ram_RW_0_r_data; // @[:anonymous source@908.4]
  wire [8:0] ram_RW_0_r_addr; // @[:anonymous source@908.4]
  wire [63:0] ram_RW_0_w_data; // @[:anonymous source@908.4]
  wire [8:0] ram_RW_0_w_addr; // @[:anonymous source@908.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@908.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@908.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [8:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@908.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = 1'h1;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@920.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@908.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_hi_us_ext( // @[:anonymous source@923.2]
  input  [6:0] W0_addr, // @[:anonymous source@924.4]
  input        W0_clk, // @[:anonymous source@925.4]
  input        W0_data, // @[:anonymous source@926.4]
  input        W0_en, // @[:anonymous source@927.4]
  input        W0_mask, // @[:anonymous source@928.4]
  input  [6:0] R0_addr, // @[:anonymous source@929.4]
  input        R0_clk, // @[:anonymous source@930.4]
  output       R0_data, // @[:anonymous source@931.4]
  input        R0_en // @[:anonymous source@932.4]
);
  reg  ram [0:63]; // @[:anonymous source@934.4]
  reg [31:0] _RAND_0;
  wire  ram_R_0_data; // @[:anonymous source@934.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@934.4]
  wire  ram_W_0_data; // @[:anonymous source@934.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@934.4]
  wire  ram_W_0_mask; // @[:anonymous source@934.4]
  wire  ram_W_0_en; // @[:anonymous source@934.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@934.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@945.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@934.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_table_ext( // @[:anonymous source@952.2]
  input  [6:0]  W0_addr, // @[:anonymous source@953.4]
  input         W0_clk, // @[:anonymous source@954.4]
  input  [10:0] W0_data, // @[:anonymous source@955.4]
  input         W0_en, // @[:anonymous source@956.4]
  input         W0_mask, // @[:anonymous source@957.4]
  input  [6:0]  R0_addr, // @[:anonymous source@958.4]
  input         R0_clk, // @[:anonymous source@959.4]
  output [10:0] R0_data, // @[:anonymous source@960.4]
  input         R0_en // @[:anonymous source@961.4]
);
  reg [10:0] ram [0:63]; // @[:anonymous source@963.4]
  reg [31:0] _RAND_0;
  wire [10:0] ram_R_0_data; // @[:anonymous source@963.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@963.4]
  wire [10:0] ram_W_0_data; // @[:anonymous source@963.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@963.4]
  wire  ram_W_0_mask; // @[:anonymous source@963.4]
  wire  ram_W_0_en; // @[:anonymous source@963.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@963.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@974.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[10:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@963.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_hi_us_0_ext( // @[:anonymous source@981.2]
  input  [7:0] W0_addr, // @[:anonymous source@982.4]
  input        W0_clk, // @[:anonymous source@983.4]
  input        W0_data, // @[:anonymous source@984.4]
  input        W0_en, // @[:anonymous source@985.4]
  input        W0_mask, // @[:anonymous source@986.4]
  input  [7:0] R0_addr, // @[:anonymous source@987.4]
  input        R0_clk, // @[:anonymous source@988.4]
  output       R0_data, // @[:anonymous source@989.4]
  input        R0_en // @[:anonymous source@990.4]
);
  reg  ram [0:63]; // @[:anonymous source@992.4]
  reg [31:0] _RAND_0;
  wire  ram_R_0_data; // @[:anonymous source@992.4]
  wire [7:0] ram_R_0_addr; // @[:anonymous source@992.4]
  wire  ram_W_0_data; // @[:anonymous source@992.4]
  wire [7:0] ram_W_0_addr; // @[:anonymous source@992.4]
  wire  ram_W_0_mask; // @[:anonymous source@992.4]
  wire  ram_W_0_en; // @[:anonymous source@992.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [7:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@992.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1003.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@992.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_table_0_ext( // @[:anonymous source@1010.2]
  input  [7:0]  W0_addr, // @[:anonymous source@1011.4]
  input         W0_clk, // @[:anonymous source@1012.4]
  input  [11:0] W0_data, // @[:anonymous source@1013.4]
  input         W0_en, // @[:anonymous source@1014.4]
  input         W0_mask, // @[:anonymous source@1015.4]
  input  [7:0]  R0_addr, // @[:anonymous source@1016.4]
  input         R0_clk, // @[:anonymous source@1017.4]
  output [11:0] R0_data, // @[:anonymous source@1018.4]
  input         R0_en // @[:anonymous source@1019.4]
);
  reg [11:0] ram [0:63]; // @[:anonymous source@1021.4]
  reg [31:0] _RAND_0;
  wire [11:0] ram_R_0_data; // @[:anonymous source@1021.4]
  wire [7:0] ram_R_0_addr; // @[:anonymous source@1021.4]
  wire [11:0] ram_W_0_data; // @[:anonymous source@1021.4]
  wire [7:0] ram_W_0_addr; // @[:anonymous source@1021.4]
  wire  ram_W_0_mask; // @[:anonymous source@1021.4]
  wire  ram_W_0_en; // @[:anonymous source@1021.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [7:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1021.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1032.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[11:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1021.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_table_1_ext( // @[:anonymous source@1039.2]
  input  [6:0]  W0_addr, // @[:anonymous source@1040.4]
  input         W0_clk, // @[:anonymous source@1041.4]
  input  [12:0] W0_data, // @[:anonymous source@1042.4]
  input         W0_en, // @[:anonymous source@1043.4]
  input         W0_mask, // @[:anonymous source@1044.4]
  input  [6:0]  R0_addr, // @[:anonymous source@1045.4]
  input         R0_clk, // @[:anonymous source@1046.4]
  output [12:0] R0_data, // @[:anonymous source@1047.4]
  input         R0_en // @[:anonymous source@1048.4]
);
  reg [12:0] ram [0:63]; // @[:anonymous source@1050.4]
  reg [31:0] _RAND_0;
  wire [12:0] ram_R_0_data; // @[:anonymous source@1050.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@1050.4]
  wire [12:0] ram_W_0_data; // @[:anonymous source@1050.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@1050.4]
  wire  ram_W_0_mask; // @[:anonymous source@1050.4]
  wire  ram_W_0_en; // @[:anonymous source@1050.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1050.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1061.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[12:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1050.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_meta_0_ext( // @[:anonymous source@1068.2]
  input  [6:0]  W0_addr, // @[:anonymous source@1069.4]
  input         W0_clk, // @[:anonymous source@1070.4]
  input  [30:0] W0_data, // @[:anonymous source@1071.4]
  input         W0_en, // @[:anonymous source@1072.4]
  input         W0_mask, // @[:anonymous source@1073.4]
  input  [6:0]  R0_addr, // @[:anonymous source@1074.4]
  input         R0_clk, // @[:anonymous source@1075.4]
  output [30:0] R0_data, // @[:anonymous source@1076.4]
  input         R0_en // @[:anonymous source@1077.4]
);
  reg [30:0] ram [0:63]; // @[:anonymous source@1079.4]
  reg [31:0] _RAND_0;
  wire [30:0] ram_R_0_data; // @[:anonymous source@1079.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@1079.4]
  wire [30:0] ram_W_0_data; // @[:anonymous source@1079.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@1079.4]
  wire  ram_W_0_mask; // @[:anonymous source@1079.4]
  wire  ram_W_0_en; // @[:anonymous source@1079.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1079.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1090.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[30:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1079.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_btb_0_ext( // @[:anonymous source@1097.2]
  input  [6:0]  W0_addr, // @[:anonymous source@1098.4]
  input         W0_clk, // @[:anonymous source@1099.4]
  input  [13:0] W0_data, // @[:anonymous source@1100.4]
  input         W0_en, // @[:anonymous source@1101.4]
  input         W0_mask, // @[:anonymous source@1102.4]
  input  [6:0]  R0_addr, // @[:anonymous source@1103.4]
  input         R0_clk, // @[:anonymous source@1104.4]
  output [13:0] R0_data, // @[:anonymous source@1105.4]
  input         R0_en // @[:anonymous source@1106.4]
);
  reg [13:0] ram [0:63]; // @[:anonymous source@1108.4]
  reg [31:0] _RAND_0;
  wire [13:0] ram_R_0_data; // @[:anonymous source@1108.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@1108.4]
  wire [13:0] ram_W_0_data; // @[:anonymous source@1108.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@1108.4]
  wire  ram_W_0_mask; // @[:anonymous source@1108.4]
  wire  ram_W_0_en; // @[:anonymous source@1108.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1108.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1119.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[13:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1108.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_ebtb_ext( // @[:anonymous source@1126.2]
  input  [6:0]  W0_addr, // @[:anonymous source@1127.4]
  input         W0_clk, // @[:anonymous source@1128.4]
  input  [39:0] W0_data, // @[:anonymous source@1129.4]
  input         W0_en, // @[:anonymous source@1130.4]
  input  [6:0]  R0_addr, // @[:anonymous source@1131.4]
  input         R0_clk, // @[:anonymous source@1132.4]
  output [39:0] R0_data, // @[:anonymous source@1133.4]
  input         R0_en // @[:anonymous source@1134.4]
);
  reg [39:0] ram [0:63]; // @[:anonymous source@1136.4]
  reg [63:0] _RAND_0;
  wire [39:0] ram_R_0_data; // @[:anonymous source@1136.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@1136.4]
  wire [39:0] ram_W_0_data; // @[:anonymous source@1136.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@1136.4]
  wire  ram_W_0_mask; // @[:anonymous source@1136.4]
  wire  ram_W_0_en; // @[:anonymous source@1136.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1136.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = 1'h1;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1147.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[39:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1136.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_data_ext( // @[:anonymous source@1154.2]
  input  [10:0] W0_addr, // @[:anonymous source@1155.4]
  input         W0_clk, // @[:anonymous source@1156.4]
  input  [1:0]  W0_data, // @[:anonymous source@1157.4]
  input         W0_en, // @[:anonymous source@1158.4]
  input         W0_mask, // @[:anonymous source@1159.4]
  input  [10:0] R0_addr, // @[:anonymous source@1160.4]
  input         R0_clk, // @[:anonymous source@1161.4]
  output [1:0]  R0_data, // @[:anonymous source@1162.4]
  input         R0_en // @[:anonymous source@1163.4]
);
  reg [1:0] ram [0:63]; // @[:anonymous source@1165.4]
  reg [31:0] _RAND_0;
  wire [1:0] ram_R_0_data; // @[:anonymous source@1165.4]
  wire [10:0] ram_R_0_addr; // @[:anonymous source@1165.4]
  wire [1:0] ram_W_0_data; // @[:anonymous source@1165.4]
  wire [10:0] ram_W_0_addr; // @[:anonymous source@1165.4]
  wire  ram_W_0_mask; // @[:anonymous source@1165.4]
  wire  ram_W_0_en; // @[:anonymous source@1165.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [10:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1165.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1176.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    ram[initvar] = _RAND_0[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[10:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1165.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_meta_ext( // @[:anonymous source@1183.2]
  input  [4:0]   W0_addr, // @[:anonymous source@1184.4]
  input          W0_clk, // @[:anonymous source@1185.4]
  input  [119:0] W0_data, // @[:anonymous source@1186.4]
  input          W0_en, // @[:anonymous source@1187.4]
  input  [4:0]   R0_addr, // @[:anonymous source@1188.4]
  input          R0_clk, // @[:anonymous source@1189.4]
  output [119:0] R0_data, // @[:anonymous source@1190.4]
  input          R0_en // @[:anonymous source@1191.4]
);
  reg [119:0] ram [0:31]; // @[:anonymous source@1193.4]
  reg [127:0] _RAND_0;
  wire [119:0] ram_R_0_data; // @[:anonymous source@1193.4]
  wire [4:0] ram_R_0_addr; // @[:anonymous source@1193.4]
  wire [119:0] ram_W_0_data; // @[:anonymous source@1193.4]
  wire [4:0] ram_W_0_addr; // @[:anonymous source@1193.4]
  wire  ram_W_0_mask; // @[:anonymous source@1193.4]
  wire  ram_W_0_en; // @[:anonymous source@1193.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [4:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1193.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = 1'h1;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1204.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram[initvar] = _RAND_0[119:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1193.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_ghist_0_ext( // @[:anonymous source@1211.2]
  input  [4:0]  W0_addr, // @[:anonymous source@1212.4]
  input         W0_clk, // @[:anonymous source@1213.4]
  input  [71:0] W0_data, // @[:anonymous source@1214.4]
  input         W0_en, // @[:anonymous source@1215.4]
  input  [4:0]  R0_addr, // @[:anonymous source@1216.4]
  input         R0_clk, // @[:anonymous source@1217.4]
  output [71:0] R0_data, // @[:anonymous source@1218.4]
  input         R0_en // @[:anonymous source@1219.4]
);
  reg [71:0] ram [0:31]; // @[:anonymous source@1221.4]
  reg [95:0] _RAND_0;
  wire [71:0] ram_R_0_data; // @[:anonymous source@1221.4]
  wire [4:0] ram_R_0_addr; // @[:anonymous source@1221.4]
  wire [71:0] ram_W_0_data; // @[:anonymous source@1221.4]
  wire [4:0] ram_W_0_addr; // @[:anonymous source@1221.4]
  wire  ram_W_0_mask; // @[:anonymous source@1221.4]
  wire  ram_W_0_en; // @[:anonymous source@1221.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [4:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1221.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = 1'h1;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1232.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {3{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram[initvar] = _RAND_0[71:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1221.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_rob_debug_inst_mem_ext( // @[:anonymous source@1239.2]
  input  [4:0]  W0_addr, // @[:anonymous source@1240.4]
  input         W0_clk, // @[:anonymous source@1241.4]
  input  [31:0] W0_data, // @[:anonymous source@1242.4]
  input         W0_en, // @[:anonymous source@1243.4]
  input         W0_mask, // @[:anonymous source@1244.4]
  input  [4:0]  R0_addr, // @[:anonymous source@1245.4]
  input         R0_clk, // @[:anonymous source@1246.4]
  output [31:0] R0_data, // @[:anonymous source@1247.4]
  input         R0_en // @[:anonymous source@1248.4]
);
  reg [31:0] ram [0:31]; // @[:anonymous source@1250.4]
  reg [31:0] _RAND_0;
  wire [31:0] ram_R_0_data; // @[:anonymous source@1250.4]
  wire [4:0] ram_R_0_addr; // @[:anonymous source@1250.4]
  wire [31:0] ram_W_0_data; // @[:anonymous source@1250.4]
  wire [4:0] ram_W_0_addr; // @[:anonymous source@1250.4]
  wire  ram_W_0_mask; // @[:anonymous source@1250.4]
  wire  ram_W_0_en; // @[:anonymous source@1250.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [4:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1250.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1261.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1250.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_l2_tlb_ram_ext( // @[:anonymous source@1268.2]
  input  [9:0]  RW0_addr, // @[:anonymous source@1269.4]
  input         RW0_clk, // @[:anonymous source@1270.4]
  input  [43:0] RW0_wdata, // @[:anonymous source@1271.4]
  output [43:0] RW0_rdata, // @[:anonymous source@1272.4]
  input         RW0_en, // @[:anonymous source@1273.4]
  input         RW0_wmode // @[:anonymous source@1274.4]
);
  reg [43:0] ram [0:63]; // @[:anonymous source@1276.4]
  reg [63:0] _RAND_0;
  wire [43:0] ram_RW_0_r_data; // @[:anonymous source@1276.4]
  wire [9:0] ram_RW_0_r_addr; // @[:anonymous source@1276.4]
  wire [43:0] ram_RW_0_w_data; // @[:anonymous source@1276.4]
  wire [9:0] ram_RW_0_w_addr; // @[:anonymous source@1276.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@1276.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@1276.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [9:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@1276.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = 1'h1;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@1288.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    ram[initvar] = _RAND_0[43:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@1276.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
